/////////////////////////////////////////////////////////////////////////////////////
// File Name : yapp.svh
// Version   : 0.1
//-------------------yapp.svh------------------------------------
/////////////////////////////////////////////////////////////////////////////////////

    
`ifndef YAPP_SVH
`define YAPP_SVH
  typedef uvm_config_db#(virtual yapp_if) yapp_vif_config;
  `include "yapp_packet.sv"
  `include "yapp_tx_monitor.sv"
  `include "yapp_tx_sequencer.sv"	
  `include "yapp_tx_seqs.sv"
  `include "yapp_tx_driver.sv"
  `include "yapp_tx_agent.sv"
  `include "yapp_env.sv"
  `include "../channel/sv/channel.svh"
  `include "router_tb.sv"

`endif// YAPP_SVH


