/////////////////////////////////////////////////////////////////////////////////////
// File Name : yapp.svh
// Version   : 0.1
//-------------------yapp.svh------------------------------------
/////////////////////////////////////////////////////////////////////////////////////

    
`ifndef YAPP_SVH
`define YAPP_SVH

  `include "yapp_packet.sv"
  `include "yapp_tx_monitor.sv"
  `include "yapp_tx_sequencer.sv"	
  `include "yapp_tx_seqs.sv"
  `include "yapp_tx_driver.sv"
  `include "yapp_tx_agent.sv"
  `include "yapp_env.sv"

`endif// YAPP_SVH


