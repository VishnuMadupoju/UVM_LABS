////////////////////////////////////////////////////////////////////////////////////////////////
// File Name : yapp_tx_seqs.sv
// version   : 0.1
// -------------yapp_tx_seqs---------------------------------------
/////////////////////////////////////////////////////////////////////////////////////////////////
